// CST455_Midterm.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module CST455_Midterm (
		input  wire        clk_clk,            //         clk.clk
		output wire [6:0]  hex0_export,        //        hex0.export
		output wire [6:0]  hex1_export,        //        hex1.export
		output wire [6:0]  hex2_export,        //        hex2.export
		output wire [6:0]  hex3_export,        //        hex3.export
		output wire [6:0]  hex4_export,        //        hex4.export
		output wire [6:0]  hex5_export,        //        hex5.export
		output wire [9:0]  leds_export,        //        leds.export
		input  wire [3:0]  pushbuttons_export, // pushbuttons.export
		output wire        sdram_clk_clk,      //   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,    //  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,      //            .ba
		output wire        sdram_wire_cas_n,   //            .cas_n
		output wire        sdram_wire_cke,     //            .cke
		output wire        sdram_wire_cs_n,    //            .cs_n
		inout  wire [15:0] sdram_wire_dq,      //            .dq
		output wire [1:0]  sdram_wire_dqm,     //            .dqm
		output wire        sdram_wire_ras_n,   //            .ras_n
		output wire        sdram_wire_we_n,    //            .we_n
		input  wire [9:0]  sw_export           //          sw.export
	);

	wire         clocks_sys_clk_clk;                                            // CLOCKS:sys_clk_clk -> [CST455_Midterm:clk, DEBUG:clk, LEDs_0:clk, Pushbuttons_0:clk, SDRAM:clk, SevenSegDecoder_0:clk, SevenSegDecoder_1:clk, SevenSegDecoder_2:clk, SevenSegDecoder_3:clk, SevenSegDecoder_4:clk, SevenSegDecoder_5:clk, Switches_0:clk, irq_mapper:clk, mm_interconnect_0:CLOCKS_sys_clk_clk, rst_controller:clk, sys_clk:clk]
	wire         cst455_midterm_debug_reset_request_reset;                      // CST455_Midterm:debug_reset_request -> [CLOCKS:ref_reset_reset, rst_controller:reset_in0]
	wire  [31:0] cst455_midterm_data_master_readdata;                           // mm_interconnect_0:CST455_Midterm_data_master_readdata -> CST455_Midterm:d_readdata
	wire         cst455_midterm_data_master_waitrequest;                        // mm_interconnect_0:CST455_Midterm_data_master_waitrequest -> CST455_Midterm:d_waitrequest
	wire         cst455_midterm_data_master_debugaccess;                        // CST455_Midterm:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CST455_Midterm_data_master_debugaccess
	wire  [27:0] cst455_midterm_data_master_address;                            // CST455_Midterm:d_address -> mm_interconnect_0:CST455_Midterm_data_master_address
	wire   [3:0] cst455_midterm_data_master_byteenable;                         // CST455_Midterm:d_byteenable -> mm_interconnect_0:CST455_Midterm_data_master_byteenable
	wire         cst455_midterm_data_master_read;                               // CST455_Midterm:d_read -> mm_interconnect_0:CST455_Midterm_data_master_read
	wire         cst455_midterm_data_master_write;                              // CST455_Midterm:d_write -> mm_interconnect_0:CST455_Midterm_data_master_write
	wire  [31:0] cst455_midterm_data_master_writedata;                          // CST455_Midterm:d_writedata -> mm_interconnect_0:CST455_Midterm_data_master_writedata
	wire  [31:0] cst455_midterm_instruction_master_readdata;                    // mm_interconnect_0:CST455_Midterm_instruction_master_readdata -> CST455_Midterm:i_readdata
	wire         cst455_midterm_instruction_master_waitrequest;                 // mm_interconnect_0:CST455_Midterm_instruction_master_waitrequest -> CST455_Midterm:i_waitrequest
	wire  [27:0] cst455_midterm_instruction_master_address;                     // CST455_Midterm:i_address -> mm_interconnect_0:CST455_Midterm_instruction_master_address
	wire         cst455_midterm_instruction_master_read;                        // CST455_Midterm:i_read -> mm_interconnect_0:CST455_Midterm_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;          // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;            // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;         // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;             // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;                // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;               // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;           // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire         mm_interconnect_0_leds_0_avalon_slave_0_chipselect;            // mm_interconnect_0:LEDs_0_avalon_slave_0_chipselect -> LEDs_0:chipselect
	wire  [31:0] mm_interconnect_0_leds_0_avalon_slave_0_readdata;              // LEDs_0:readdata -> mm_interconnect_0:LEDs_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_leds_0_avalon_slave_0_address;               // mm_interconnect_0:LEDs_0_avalon_slave_0_address -> LEDs_0:address
	wire         mm_interconnect_0_leds_0_avalon_slave_0_read;                  // mm_interconnect_0:LEDs_0_avalon_slave_0_read -> LEDs_0:read
	wire         mm_interconnect_0_leds_0_avalon_slave_0_write;                 // mm_interconnect_0:LEDs_0_avalon_slave_0_write -> LEDs_0:write
	wire  [31:0] mm_interconnect_0_leds_0_avalon_slave_0_writedata;             // mm_interconnect_0:LEDs_0_avalon_slave_0_writedata -> LEDs_0:writedata
	wire         mm_interconnect_0_switches_0_avalon_slave_0_chipselect;        // mm_interconnect_0:Switches_0_avalon_slave_0_chipselect -> Switches_0:chipselect
	wire  [31:0] mm_interconnect_0_switches_0_avalon_slave_0_readdata;          // Switches_0:readdata -> mm_interconnect_0:Switches_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_switches_0_avalon_slave_0_address;           // mm_interconnect_0:Switches_0_avalon_slave_0_address -> Switches_0:address
	wire         mm_interconnect_0_switches_0_avalon_slave_0_read;              // mm_interconnect_0:Switches_0_avalon_slave_0_read -> Switches_0:read
	wire         mm_interconnect_0_pushbuttons_0_avalon_slave_0_chipselect;     // mm_interconnect_0:Pushbuttons_0_avalon_slave_0_chipselect -> Pushbuttons_0:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_0_avalon_slave_0_readdata;       // Pushbuttons_0:readdata -> mm_interconnect_0:Pushbuttons_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_0_avalon_slave_0_address;        // mm_interconnect_0:Pushbuttons_0_avalon_slave_0_address -> Pushbuttons_0:address
	wire         mm_interconnect_0_pushbuttons_0_avalon_slave_0_read;           // mm_interconnect_0:Pushbuttons_0_avalon_slave_0_read -> Pushbuttons_0:read
	wire         mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_chipselect -> SevenSegDecoder_1:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_readdata;   // SevenSegDecoder_1:readdata -> mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_address -> SevenSegDecoder_1:address
	wire         mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_write -> SevenSegDecoder_1:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_writedata -> SevenSegDecoder_1:writedata
	wire         mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_chipselect -> SevenSegDecoder_2:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_readdata;   // SevenSegDecoder_2:readdata -> mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_address -> SevenSegDecoder_2:address
	wire         mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_write -> SevenSegDecoder_2:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_writedata -> SevenSegDecoder_2:writedata
	wire         mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_chipselect -> SevenSegDecoder_4:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_readdata;   // SevenSegDecoder_4:readdata -> mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_address -> SevenSegDecoder_4:address
	wire         mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_write -> SevenSegDecoder_4:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_writedata -> SevenSegDecoder_4:writedata
	wire         mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_chipselect -> SevenSegDecoder_5:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_readdata;   // SevenSegDecoder_5:readdata -> mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_address -> SevenSegDecoder_5:address
	wire         mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_write -> SevenSegDecoder_5:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_writedata -> SevenSegDecoder_5:writedata
	wire         mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_chipselect -> SevenSegDecoder_3:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_readdata;   // SevenSegDecoder_3:readdata -> mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_address -> SevenSegDecoder_3:address
	wire         mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_write -> SevenSegDecoder_3:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_writedata -> SevenSegDecoder_3:writedata
	wire         mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_chipselect -> SevenSegDecoder_0:chipselect
	wire  [31:0] mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_readdata;   // SevenSegDecoder_0:readdata -> mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_address -> SevenSegDecoder_0:address
	wire         mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_write -> SevenSegDecoder_0:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_writedata -> SevenSegDecoder_0:writedata
	wire  [31:0] mm_interconnect_0_cst455_midterm_debug_mem_slave_readdata;     // CST455_Midterm:debug_mem_slave_readdata -> mm_interconnect_0:CST455_Midterm_debug_mem_slave_readdata
	wire         mm_interconnect_0_cst455_midterm_debug_mem_slave_waitrequest;  // CST455_Midterm:debug_mem_slave_waitrequest -> mm_interconnect_0:CST455_Midterm_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cst455_midterm_debug_mem_slave_debugaccess;  // mm_interconnect_0:CST455_Midterm_debug_mem_slave_debugaccess -> CST455_Midterm:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cst455_midterm_debug_mem_slave_address;      // mm_interconnect_0:CST455_Midterm_debug_mem_slave_address -> CST455_Midterm:debug_mem_slave_address
	wire         mm_interconnect_0_cst455_midterm_debug_mem_slave_read;         // mm_interconnect_0:CST455_Midterm_debug_mem_slave_read -> CST455_Midterm:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cst455_midterm_debug_mem_slave_byteenable;   // mm_interconnect_0:CST455_Midterm_debug_mem_slave_byteenable -> CST455_Midterm:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cst455_midterm_debug_mem_slave_write;        // mm_interconnect_0:CST455_Midterm_debug_mem_slave_write -> CST455_Midterm:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cst455_midterm_debug_mem_slave_writedata;    // mm_interconnect_0:CST455_Midterm_debug_mem_slave_writedata -> CST455_Midterm:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                         // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                           // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                        // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                            // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                               // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                         // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                      // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                              // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                          // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_sys_clk_s1_chipselect;                       // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                         // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                          // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                            // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                        // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         irq_mapper_receiver0_irq;                                      // sys_clk:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // DEBUG:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cst455_midterm_irq_irq;                                        // irq_mapper:sender_irq -> CST455_Midterm:irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [CST455_Midterm:reset_n, DEBUG:rst_n, LEDs_0:reset_n, Pushbuttons_0:reset_n, SDRAM:reset_n, SevenSegDecoder_0:reset_n, SevenSegDecoder_1:reset_n, SevenSegDecoder_2:reset_n, SevenSegDecoder_3:reset_n, SevenSegDecoder_4:reset_n, SevenSegDecoder_5:reset_n, Switches_0:reset_n, irq_mapper:reset, mm_interconnect_0:CST455_Midterm_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sys_clk:reset_n]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [CST455_Midterm:reset_req, rst_translator:reset_req_in]

	CST455_Midterm_CLOCKS clocks (
		.ref_clk_clk        (clk_clk),                                  //      ref_clk.clk
		.ref_reset_reset    (cst455_midterm_debug_reset_request_reset), //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),                       //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                            //    sdram_clk.clk
		.reset_source_reset ()                                          // reset_source.reset
	);

	CST455_Midterm_CST455_Midterm cst455_midterm (
		.clk                                 (clocks_sys_clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                              //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                           (cst455_midterm_data_master_address),                           //               data_master.address
		.d_byteenable                        (cst455_midterm_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cst455_midterm_data_master_read),                              //                          .read
		.d_readdata                          (cst455_midterm_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cst455_midterm_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cst455_midterm_data_master_write),                             //                          .write
		.d_writedata                         (cst455_midterm_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cst455_midterm_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cst455_midterm_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cst455_midterm_instruction_master_read),                       //                          .read
		.i_readdata                          (cst455_midterm_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cst455_midterm_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cst455_midterm_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cst455_midterm_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cst455_midterm_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cst455_midterm_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cst455_midterm_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cst455_midterm_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cst455_midterm_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cst455_midterm_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cst455_midterm_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cst455_midterm_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                              // custom_instruction_master.readra
	);

	CST455_Midterm_DEBUG debug (
		.clk            (clocks_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                               //               irq.irq
	);

	LEDController leds_0 (
		.address    (mm_interconnect_0_leds_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_leds_0_avalon_slave_0_chipselect), //               .chipselect
		.read       (mm_interconnect_0_leds_0_avalon_slave_0_read),       //               .read
		.write      (mm_interconnect_0_leds_0_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_leds_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_leds_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clocks_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //          reset.reset_n
		.led_out    (leds_export)                                         //    conduit_end.export
	);

	PushbuttonReader pushbuttons_0 (
		.address     (mm_interconnect_0_pushbuttons_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect  (mm_interconnect_0_pushbuttons_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata    (mm_interconnect_0_pushbuttons_0_avalon_slave_0_readdata),   //               .readdata
		.read        (mm_interconnect_0_pushbuttons_0_avalon_slave_0_read),       //               .read
		.clk         (clocks_sys_clk_clk),                                        //          clock.clk
		.reset_n     (~rst_controller_reset_out_reset),                           //          reset.reset_n
		.pushbuttons (pushbuttons_export)                                         //    conduit_end.export
	);

	CST455_Midterm_SDRAM sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	SevenSegDecoder sevensegdecoder_0 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex0_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_1 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex1_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_2 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex2_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_3 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex3_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_4 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex4_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_5 (
		.clk        (clocks_sys_clk_clk),                                            //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_readdata),   //               .readdata
		.segs       (hex5_export)                                                    //    conduit_end.export
	);

	SwitchReader switches_0 (
		.address    (mm_interconnect_0_switches_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_switches_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_switches_0_avalon_slave_0_readdata),   //               .readdata
		.read       (mm_interconnect_0_switches_0_avalon_slave_0_read),       //               .read
		.clk        (clocks_sys_clk_clk),                                     //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //          reset.reset_n
		.switch     (sw_export)                                               //    conduit_end.export
	);

	CST455_Midterm_sys_clk sys_clk (
		.clk        (clocks_sys_clk_clk),                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	CST455_Midterm_mm_interconnect_0 mm_interconnect_0 (
		.CLOCKS_sys_clk_clk                               (clocks_sys_clk_clk),                                            //                             CLOCKS_sys_clk.clk
		.CST455_Midterm_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // CST455_Midterm_reset_reset_bridge_in_reset.reset
		.CST455_Midterm_data_master_address               (cst455_midterm_data_master_address),                            //                 CST455_Midterm_data_master.address
		.CST455_Midterm_data_master_waitrequest           (cst455_midterm_data_master_waitrequest),                        //                                           .waitrequest
		.CST455_Midterm_data_master_byteenable            (cst455_midterm_data_master_byteenable),                         //                                           .byteenable
		.CST455_Midterm_data_master_read                  (cst455_midterm_data_master_read),                               //                                           .read
		.CST455_Midterm_data_master_readdata              (cst455_midterm_data_master_readdata),                           //                                           .readdata
		.CST455_Midterm_data_master_write                 (cst455_midterm_data_master_write),                              //                                           .write
		.CST455_Midterm_data_master_writedata             (cst455_midterm_data_master_writedata),                          //                                           .writedata
		.CST455_Midterm_data_master_debugaccess           (cst455_midterm_data_master_debugaccess),                        //                                           .debugaccess
		.CST455_Midterm_instruction_master_address        (cst455_midterm_instruction_master_address),                     //          CST455_Midterm_instruction_master.address
		.CST455_Midterm_instruction_master_waitrequest    (cst455_midterm_instruction_master_waitrequest),                 //                                           .waitrequest
		.CST455_Midterm_instruction_master_read           (cst455_midterm_instruction_master_read),                        //                                           .read
		.CST455_Midterm_instruction_master_readdata       (cst455_midterm_instruction_master_readdata),                    //                                           .readdata
		.CST455_Midterm_debug_mem_slave_address           (mm_interconnect_0_cst455_midterm_debug_mem_slave_address),      //             CST455_Midterm_debug_mem_slave.address
		.CST455_Midterm_debug_mem_slave_write             (mm_interconnect_0_cst455_midterm_debug_mem_slave_write),        //                                           .write
		.CST455_Midterm_debug_mem_slave_read              (mm_interconnect_0_cst455_midterm_debug_mem_slave_read),         //                                           .read
		.CST455_Midterm_debug_mem_slave_readdata          (mm_interconnect_0_cst455_midterm_debug_mem_slave_readdata),     //                                           .readdata
		.CST455_Midterm_debug_mem_slave_writedata         (mm_interconnect_0_cst455_midterm_debug_mem_slave_writedata),    //                                           .writedata
		.CST455_Midterm_debug_mem_slave_byteenable        (mm_interconnect_0_cst455_midterm_debug_mem_slave_byteenable),   //                                           .byteenable
		.CST455_Midterm_debug_mem_slave_waitrequest       (mm_interconnect_0_cst455_midterm_debug_mem_slave_waitrequest),  //                                           .waitrequest
		.CST455_Midterm_debug_mem_slave_debugaccess       (mm_interconnect_0_cst455_midterm_debug_mem_slave_debugaccess),  //                                           .debugaccess
		.DEBUG_avalon_jtag_slave_address                  (mm_interconnect_0_debug_avalon_jtag_slave_address),             //                    DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write                    (mm_interconnect_0_debug_avalon_jtag_slave_write),               //                                           .write
		.DEBUG_avalon_jtag_slave_read                     (mm_interconnect_0_debug_avalon_jtag_slave_read),                //                                           .read
		.DEBUG_avalon_jtag_slave_readdata                 (mm_interconnect_0_debug_avalon_jtag_slave_readdata),            //                                           .readdata
		.DEBUG_avalon_jtag_slave_writedata                (mm_interconnect_0_debug_avalon_jtag_slave_writedata),           //                                           .writedata
		.DEBUG_avalon_jtag_slave_waitrequest              (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),         //                                           .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect               (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),          //                                           .chipselect
		.LEDs_0_avalon_slave_0_address                    (mm_interconnect_0_leds_0_avalon_slave_0_address),               //                      LEDs_0_avalon_slave_0.address
		.LEDs_0_avalon_slave_0_write                      (mm_interconnect_0_leds_0_avalon_slave_0_write),                 //                                           .write
		.LEDs_0_avalon_slave_0_read                       (mm_interconnect_0_leds_0_avalon_slave_0_read),                  //                                           .read
		.LEDs_0_avalon_slave_0_readdata                   (mm_interconnect_0_leds_0_avalon_slave_0_readdata),              //                                           .readdata
		.LEDs_0_avalon_slave_0_writedata                  (mm_interconnect_0_leds_0_avalon_slave_0_writedata),             //                                           .writedata
		.LEDs_0_avalon_slave_0_chipselect                 (mm_interconnect_0_leds_0_avalon_slave_0_chipselect),            //                                           .chipselect
		.Pushbuttons_0_avalon_slave_0_address             (mm_interconnect_0_pushbuttons_0_avalon_slave_0_address),        //               Pushbuttons_0_avalon_slave_0.address
		.Pushbuttons_0_avalon_slave_0_read                (mm_interconnect_0_pushbuttons_0_avalon_slave_0_read),           //                                           .read
		.Pushbuttons_0_avalon_slave_0_readdata            (mm_interconnect_0_pushbuttons_0_avalon_slave_0_readdata),       //                                           .readdata
		.Pushbuttons_0_avalon_slave_0_chipselect          (mm_interconnect_0_pushbuttons_0_avalon_slave_0_chipselect),     //                                           .chipselect
		.SDRAM_s1_address                                 (mm_interconnect_0_sdram_s1_address),                            //                                   SDRAM_s1.address
		.SDRAM_s1_write                                   (mm_interconnect_0_sdram_s1_write),                              //                                           .write
		.SDRAM_s1_read                                    (mm_interconnect_0_sdram_s1_read),                               //                                           .read
		.SDRAM_s1_readdata                                (mm_interconnect_0_sdram_s1_readdata),                           //                                           .readdata
		.SDRAM_s1_writedata                               (mm_interconnect_0_sdram_s1_writedata),                          //                                           .writedata
		.SDRAM_s1_byteenable                              (mm_interconnect_0_sdram_s1_byteenable),                         //                                           .byteenable
		.SDRAM_s1_readdatavalid                           (mm_interconnect_0_sdram_s1_readdatavalid),                      //                                           .readdatavalid
		.SDRAM_s1_waitrequest                             (mm_interconnect_0_sdram_s1_waitrequest),                        //                                           .waitrequest
		.SDRAM_s1_chipselect                              (mm_interconnect_0_sdram_s1_chipselect),                         //                                           .chipselect
		.SevenSegDecoder_0_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address),    //           SevenSegDecoder_0_avalon_slave_0.address
		.SevenSegDecoder_0_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_0_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_0_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_0_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect), //                                           .chipselect
		.SevenSegDecoder_1_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address),    //           SevenSegDecoder_1_avalon_slave_0.address
		.SevenSegDecoder_1_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_1_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_1_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_1_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect), //                                           .chipselect
		.SevenSegDecoder_2_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address),    //           SevenSegDecoder_2_avalon_slave_0.address
		.SevenSegDecoder_2_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_2_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_2_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_2_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect), //                                           .chipselect
		.SevenSegDecoder_3_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address),    //           SevenSegDecoder_3_avalon_slave_0.address
		.SevenSegDecoder_3_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_3_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_3_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_3_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect), //                                           .chipselect
		.SevenSegDecoder_4_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address),    //           SevenSegDecoder_4_avalon_slave_0.address
		.SevenSegDecoder_4_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_4_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_4_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_4_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect), //                                           .chipselect
		.SevenSegDecoder_5_avalon_slave_0_address         (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address),    //           SevenSegDecoder_5_avalon_slave_0.address
		.SevenSegDecoder_5_avalon_slave_0_write           (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write),      //                                           .write
		.SevenSegDecoder_5_avalon_slave_0_readdata        (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_readdata),   //                                           .readdata
		.SevenSegDecoder_5_avalon_slave_0_writedata       (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata),  //                                           .writedata
		.SevenSegDecoder_5_avalon_slave_0_chipselect      (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect), //                                           .chipselect
		.Switches_0_avalon_slave_0_address                (mm_interconnect_0_switches_0_avalon_slave_0_address),           //                  Switches_0_avalon_slave_0.address
		.Switches_0_avalon_slave_0_read                   (mm_interconnect_0_switches_0_avalon_slave_0_read),              //                                           .read
		.Switches_0_avalon_slave_0_readdata               (mm_interconnect_0_switches_0_avalon_slave_0_readdata),          //                                           .readdata
		.Switches_0_avalon_slave_0_chipselect             (mm_interconnect_0_switches_0_avalon_slave_0_chipselect),        //                                           .chipselect
		.sys_clk_s1_address                               (mm_interconnect_0_sys_clk_s1_address),                          //                                 sys_clk_s1.address
		.sys_clk_s1_write                                 (mm_interconnect_0_sys_clk_s1_write),                            //                                           .write
		.sys_clk_s1_readdata                              (mm_interconnect_0_sys_clk_s1_readdata),                         //                                           .readdata
		.sys_clk_s1_writedata                             (mm_interconnect_0_sys_clk_s1_writedata),                        //                                           .writedata
		.sys_clk_s1_chipselect                            (mm_interconnect_0_sys_clk_s1_chipselect)                        //                                           .chipselect
	);

	CST455_Midterm_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cst455_midterm_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cst455_midterm_debug_reset_request_reset), // reset_in0.reset
		.clk            (clocks_sys_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_in1      (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
