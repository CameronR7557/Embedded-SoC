// Lab03.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module Lab03 (
		input  wire       clk_clk,         //      clk.clk
		output wire [6:0] hex0_export,     //     hex0.export
		output wire [6:0] hex1_export,     //     hex1.export
		output wire [6:0] hex2_export,     //     hex2.export
		input  wire [9:0] switches_export  // switches.export
	);

	wire         lab03_debug_reset_request_reset;                       // Lab03:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] lab03_data_master_readdata;                            // mm_interconnect_0:Lab03_data_master_readdata -> Lab03:d_readdata
	wire         lab03_data_master_waitrequest;                         // mm_interconnect_0:Lab03_data_master_waitrequest -> Lab03:d_waitrequest
	wire         lab03_data_master_debugaccess;                         // Lab03:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Lab03_data_master_debugaccess
	wire  [13:0] lab03_data_master_address;                             // Lab03:d_address -> mm_interconnect_0:Lab03_data_master_address
	wire   [3:0] lab03_data_master_byteenable;                          // Lab03:d_byteenable -> mm_interconnect_0:Lab03_data_master_byteenable
	wire         lab03_data_master_read;                                // Lab03:d_read -> mm_interconnect_0:Lab03_data_master_read
	wire         lab03_data_master_write;                               // Lab03:d_write -> mm_interconnect_0:Lab03_data_master_write
	wire  [31:0] lab03_data_master_writedata;                           // Lab03:d_writedata -> mm_interconnect_0:Lab03_data_master_writedata
	wire  [31:0] lab03_instruction_master_readdata;                     // mm_interconnect_0:Lab03_instruction_master_readdata -> Lab03:i_readdata
	wire         lab03_instruction_master_waitrequest;                  // mm_interconnect_0:Lab03_instruction_master_waitrequest -> Lab03:i_waitrequest
	wire  [13:0] lab03_instruction_master_address;                      // Lab03:i_address -> mm_interconnect_0:Lab03_instruction_master_address
	wire         lab03_instruction_master_read;                         // Lab03:i_read -> mm_interconnect_0:Lab03_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_lab03_debug_mem_slave_readdata;      // Lab03:debug_mem_slave_readdata -> mm_interconnect_0:Lab03_debug_mem_slave_readdata
	wire         mm_interconnect_0_lab03_debug_mem_slave_waitrequest;   // Lab03:debug_mem_slave_waitrequest -> mm_interconnect_0:Lab03_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_lab03_debug_mem_slave_debugaccess;   // mm_interconnect_0:Lab03_debug_mem_slave_debugaccess -> Lab03:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_lab03_debug_mem_slave_address;       // mm_interconnect_0:Lab03_debug_mem_slave_address -> Lab03:debug_mem_slave_address
	wire         mm_interconnect_0_lab03_debug_mem_slave_read;          // mm_interconnect_0:Lab03_debug_mem_slave_read -> Lab03:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_lab03_debug_mem_slave_byteenable;    // mm_interconnect_0:Lab03_debug_mem_slave_byteenable -> Lab03:debug_mem_slave_byteenable
	wire         mm_interconnect_0_lab03_debug_mem_slave_write;         // mm_interconnect_0:Lab03_debug_mem_slave_write -> Lab03:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_lab03_debug_mem_slave_writedata;     // mm_interconnect_0:Lab03_debug_mem_slave_writedata -> Lab03:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                  // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                    // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire   [9:0] mm_interconnect_0_sram_s1_address;                     // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                  // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                       // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                   // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                       // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_display0_s1_chipselect;              // mm_interconnect_0:DISPLAY0_s1_chipselect -> DISPLAY0:chipselect
	wire  [31:0] mm_interconnect_0_display0_s1_readdata;                // DISPLAY0:readdata -> mm_interconnect_0:DISPLAY0_s1_readdata
	wire   [2:0] mm_interconnect_0_display0_s1_address;                 // mm_interconnect_0:DISPLAY0_s1_address -> DISPLAY0:address
	wire         mm_interconnect_0_display0_s1_write;                   // mm_interconnect_0:DISPLAY0_s1_write -> DISPLAY0:write_n
	wire  [31:0] mm_interconnect_0_display0_s1_writedata;               // mm_interconnect_0:DISPLAY0_s1_writedata -> DISPLAY0:writedata
	wire         mm_interconnect_0_display1_s1_chipselect;              // mm_interconnect_0:DISPLAY1_s1_chipselect -> DISPLAY1:chipselect
	wire  [31:0] mm_interconnect_0_display1_s1_readdata;                // DISPLAY1:readdata -> mm_interconnect_0:DISPLAY1_s1_readdata
	wire   [2:0] mm_interconnect_0_display1_s1_address;                 // mm_interconnect_0:DISPLAY1_s1_address -> DISPLAY1:address
	wire         mm_interconnect_0_display1_s1_write;                   // mm_interconnect_0:DISPLAY1_s1_write -> DISPLAY1:write_n
	wire  [31:0] mm_interconnect_0_display1_s1_writedata;               // mm_interconnect_0:DISPLAY1_s1_writedata -> DISPLAY1:writedata
	wire         mm_interconnect_0_display2_s1_chipselect;              // mm_interconnect_0:DISPLAY2_s1_chipselect -> DISPLAY2:chipselect
	wire  [31:0] mm_interconnect_0_display2_s1_readdata;                // DISPLAY2:readdata -> mm_interconnect_0:DISPLAY2_s1_readdata
	wire   [2:0] mm_interconnect_0_display2_s1_address;                 // mm_interconnect_0:DISPLAY2_s1_address -> DISPLAY2:address
	wire         mm_interconnect_0_display2_s1_write;                   // mm_interconnect_0:DISPLAY2_s1_write -> DISPLAY2:write_n
	wire  [31:0] mm_interconnect_0_display2_s1_writedata;               // mm_interconnect_0:DISPLAY2_s1_writedata -> DISPLAY2:writedata
	wire         mm_interconnect_0_sw_s1_chipselect;                    // mm_interconnect_0:SW_s1_chipselect -> SW:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                      // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                       // mm_interconnect_0:SW_s1_address -> SW:address
	wire         mm_interconnect_0_sw_s1_write;                         // mm_interconnect_0:SW_s1_write -> SW:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                     // mm_interconnect_0:SW_s1_writedata -> SW:writedata
	wire         irq_mapper_receiver0_irq;                              // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] lab03_irq_irq;                                         // irq_mapper:sender_irq -> Lab03:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [DEBUG:rst_n, DISPLAY0:reset_n, DISPLAY1:reset_n, DISPLAY2:reset_n, Lab03:reset_n, SRAM:reset, SW:reset_n, irq_mapper:reset, mm_interconnect_0:Lab03_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [Lab03:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	Lab03_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	Lab03_DISPLAY0 display0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_display0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                               // external_connection.export
	);

	Lab03_DISPLAY0 display1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_display1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                               // external_connection.export
	);

	Lab03_DISPLAY0 display2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_display2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_display2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_display2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_display2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_display2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                               // external_connection.export
	);

	Lab03_Lab03 lab03 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (lab03_data_master_address),                           //               data_master.address
		.d_byteenable                        (lab03_data_master_byteenable),                        //                          .byteenable
		.d_read                              (lab03_data_master_read),                              //                          .read
		.d_readdata                          (lab03_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (lab03_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (lab03_data_master_write),                             //                          .write
		.d_writedata                         (lab03_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (lab03_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (lab03_instruction_master_address),                    //        instruction_master.address
		.i_read                              (lab03_instruction_master_read),                       //                          .read
		.i_readdata                          (lab03_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (lab03_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (lab03_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (lab03_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_lab03_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_lab03_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_lab03_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_lab03_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_lab03_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_lab03_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_lab03_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_lab03_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	Lab03_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	Lab03_SW sw (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (switches_export)                     // external_connection.export
	);

	Lab03_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                               //                         clk_0_clk.clk
		.Lab03_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // Lab03_reset_reset_bridge_in_reset.reset
		.Lab03_data_master_address               (lab03_data_master_address),                             //                 Lab03_data_master.address
		.Lab03_data_master_waitrequest           (lab03_data_master_waitrequest),                         //                                  .waitrequest
		.Lab03_data_master_byteenable            (lab03_data_master_byteenable),                          //                                  .byteenable
		.Lab03_data_master_read                  (lab03_data_master_read),                                //                                  .read
		.Lab03_data_master_readdata              (lab03_data_master_readdata),                            //                                  .readdata
		.Lab03_data_master_write                 (lab03_data_master_write),                               //                                  .write
		.Lab03_data_master_writedata             (lab03_data_master_writedata),                           //                                  .writedata
		.Lab03_data_master_debugaccess           (lab03_data_master_debugaccess),                         //                                  .debugaccess
		.Lab03_instruction_master_address        (lab03_instruction_master_address),                      //          Lab03_instruction_master.address
		.Lab03_instruction_master_waitrequest    (lab03_instruction_master_waitrequest),                  //                                  .waitrequest
		.Lab03_instruction_master_read           (lab03_instruction_master_read),                         //                                  .read
		.Lab03_instruction_master_readdata       (lab03_instruction_master_readdata),                     //                                  .readdata
		.DEBUG_avalon_jtag_slave_address         (mm_interconnect_0_debug_avalon_jtag_slave_address),     //           DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write           (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                  .write
		.DEBUG_avalon_jtag_slave_read            (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                  .read
		.DEBUG_avalon_jtag_slave_readdata        (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                  .readdata
		.DEBUG_avalon_jtag_slave_writedata       (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                  .writedata
		.DEBUG_avalon_jtag_slave_waitrequest     (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect      (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.DISPLAY0_s1_address                     (mm_interconnect_0_display0_s1_address),                 //                       DISPLAY0_s1.address
		.DISPLAY0_s1_write                       (mm_interconnect_0_display0_s1_write),                   //                                  .write
		.DISPLAY0_s1_readdata                    (mm_interconnect_0_display0_s1_readdata),                //                                  .readdata
		.DISPLAY0_s1_writedata                   (mm_interconnect_0_display0_s1_writedata),               //                                  .writedata
		.DISPLAY0_s1_chipselect                  (mm_interconnect_0_display0_s1_chipselect),              //                                  .chipselect
		.DISPLAY1_s1_address                     (mm_interconnect_0_display1_s1_address),                 //                       DISPLAY1_s1.address
		.DISPLAY1_s1_write                       (mm_interconnect_0_display1_s1_write),                   //                                  .write
		.DISPLAY1_s1_readdata                    (mm_interconnect_0_display1_s1_readdata),                //                                  .readdata
		.DISPLAY1_s1_writedata                   (mm_interconnect_0_display1_s1_writedata),               //                                  .writedata
		.DISPLAY1_s1_chipselect                  (mm_interconnect_0_display1_s1_chipselect),              //                                  .chipselect
		.DISPLAY2_s1_address                     (mm_interconnect_0_display2_s1_address),                 //                       DISPLAY2_s1.address
		.DISPLAY2_s1_write                       (mm_interconnect_0_display2_s1_write),                   //                                  .write
		.DISPLAY2_s1_readdata                    (mm_interconnect_0_display2_s1_readdata),                //                                  .readdata
		.DISPLAY2_s1_writedata                   (mm_interconnect_0_display2_s1_writedata),               //                                  .writedata
		.DISPLAY2_s1_chipselect                  (mm_interconnect_0_display2_s1_chipselect),              //                                  .chipselect
		.Lab03_debug_mem_slave_address           (mm_interconnect_0_lab03_debug_mem_slave_address),       //             Lab03_debug_mem_slave.address
		.Lab03_debug_mem_slave_write             (mm_interconnect_0_lab03_debug_mem_slave_write),         //                                  .write
		.Lab03_debug_mem_slave_read              (mm_interconnect_0_lab03_debug_mem_slave_read),          //                                  .read
		.Lab03_debug_mem_slave_readdata          (mm_interconnect_0_lab03_debug_mem_slave_readdata),      //                                  .readdata
		.Lab03_debug_mem_slave_writedata         (mm_interconnect_0_lab03_debug_mem_slave_writedata),     //                                  .writedata
		.Lab03_debug_mem_slave_byteenable        (mm_interconnect_0_lab03_debug_mem_slave_byteenable),    //                                  .byteenable
		.Lab03_debug_mem_slave_waitrequest       (mm_interconnect_0_lab03_debug_mem_slave_waitrequest),   //                                  .waitrequest
		.Lab03_debug_mem_slave_debugaccess       (mm_interconnect_0_lab03_debug_mem_slave_debugaccess),   //                                  .debugaccess
		.SRAM_s1_address                         (mm_interconnect_0_sram_s1_address),                     //                           SRAM_s1.address
		.SRAM_s1_write                           (mm_interconnect_0_sram_s1_write),                       //                                  .write
		.SRAM_s1_readdata                        (mm_interconnect_0_sram_s1_readdata),                    //                                  .readdata
		.SRAM_s1_writedata                       (mm_interconnect_0_sram_s1_writedata),                   //                                  .writedata
		.SRAM_s1_byteenable                      (mm_interconnect_0_sram_s1_byteenable),                  //                                  .byteenable
		.SRAM_s1_chipselect                      (mm_interconnect_0_sram_s1_chipselect),                  //                                  .chipselect
		.SRAM_s1_clken                           (mm_interconnect_0_sram_s1_clken),                       //                                  .clken
		.SW_s1_address                           (mm_interconnect_0_sw_s1_address),                       //                             SW_s1.address
		.SW_s1_write                             (mm_interconnect_0_sw_s1_write),                         //                                  .write
		.SW_s1_readdata                          (mm_interconnect_0_sw_s1_readdata),                      //                                  .readdata
		.SW_s1_writedata                         (mm_interconnect_0_sw_s1_writedata),                     //                                  .writedata
		.SW_s1_chipselect                        (mm_interconnect_0_sw_s1_chipselect)                     //                                  .chipselect
	);

	Lab03_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (lab03_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (lab03_debug_reset_request_reset),    // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
