//-----------------------------------------------------------------------------    
//   University: Oregon Institute of Technology – CSET Department
//   Class: CST 455
//   Author: Cameron Robinson
//   Lab: 6
//   Project: HPS and Linux
//   File Name: Lab06.v
//   List of other files used: None
//-----------------------------------------------------------------------------    
//   Sets up the connections for the DE10-Standard HPS. Instantiates the processor
//		module. Includes connections for hex0 - hex5, LED0 - LED9, and SW0 - SW9
//-----------------------------------------------------------------------------    
//   Date: 11/14/2023
//   Version: 1.0
//   Revision:
//   11/14/2023 Initial Version
//   11/15/2023 Added HEX3-5 to force all segments to turn off
//-----------------------------------------------------------------------------


//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Lab06(

	//////////// CLOCK //////////
	input 		          		CLOCK_50,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// Seg7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,		//HEX3 - HEX5 are here just to make sure all segments are turned off
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// HPS //////////
	inout 		          		HPS_CONV_USB_N,
	output		    [14:0]		HPS_DDR3_ADDR,
	output		     [2:0]		HPS_DDR3_BA,
	output		          		HPS_DDR3_CAS_N,
	output		          		HPS_DDR3_CKE,
	output		          		HPS_DDR3_CK_N,
	output		          		HPS_DDR3_CK_P,
	output		          		HPS_DDR3_CS_N,
	output		     [3:0]		HPS_DDR3_DM,
	inout 		    [31:0]		HPS_DDR3_DQ,
	inout 		     [3:0]		HPS_DDR3_DQS_N,
	inout 		     [3:0]		HPS_DDR3_DQS_P,
	output		          		HPS_DDR3_ODT,
	output		          		HPS_DDR3_RAS_N,
	output		          		HPS_DDR3_RESET_N,
	input 		          		HPS_DDR3_RZQ,
	output		          		HPS_DDR3_WE_N,
	output		          		HPS_ENET_GTX_CLK,
	inout 		          		HPS_ENET_INT_N,
	output		          		HPS_ENET_MDC,
	inout 		          		HPS_ENET_MDIO,
	input 		          		HPS_ENET_RX_CLK,
	input 		     [3:0]		HPS_ENET_RX_DATA,
	input 		          		HPS_ENET_RX_DV,
	output		     [3:0]		HPS_ENET_TX_DATA,
	output		          		HPS_ENET_TX_EN,
	inout 		     [3:0]		HPS_FLASH_DATA,
	output		          		HPS_FLASH_DCLK,
	output		          		HPS_FLASH_NCSO,
	inout 		          		HPS_GSENSOR_INT,
	inout 		          		HPS_I2C1_SCLK,
	inout 		          		HPS_I2C1_SDAT,
	inout 		          		HPS_I2C2_SCLK,
	inout 		          		HPS_I2C2_SDAT,
	inout 		          		HPS_I2C_CONTROL,
	inout 		          		HPS_KEY,
	inout 		          		HPS_LCM_BK,
	inout 		          		HPS_LCM_D_C,
	inout 		          		HPS_LCM_RST_N,
	output		          		HPS_LCM_SPIM_CLK,
	input 		          		HPS_LCM_SPIM_MISO,
	output		          		HPS_LCM_SPIM_MOSI,
	output		          		HPS_LCM_SPIM_SS,
	inout 		          		HPS_LED,
	inout 		          		HPS_LTC_GPIO,
	output		          		HPS_SD_CLK,
	inout 		          		HPS_SD_CMD,
	inout 		     [3:0]		HPS_SD_DATA,
	output		          		HPS_SPIM_CLK,
	input 		          		HPS_SPIM_MISO,
	output		          		HPS_SPIM_MOSI,
	output		          		HPS_SPIM_SS,
	input 		          		HPS_UART_RX,
	output		          		HPS_UART_TX,
	input 		          		HPS_USB_CLKOUT,
	inout 		     [7:0]		HPS_USB_DATA,
	input 		          		HPS_USB_DIR,
	input 		          		HPS_USB_NXT,
	output		          		HPS_USB_STP
);



//=======================================================
//  REG/WIRE declarations
//=======================================================




//=======================================================
//  Structural coding
//=======================================================
	 
    Lab06_HPS u0 (
        .clk_clk                         (CLOCK_50),                    //         clk.clk
        .hex0_export                     (HEX0),                     	//     	  hex0.export
        .hex1_export                     (HEX1),                     	//         hex1.export
        .hex2_export                     (HEX2),                     	//         hex2.export
        .hps_io_hps_io_emac1_inst_TX_CLK (HPS_ENET_GTX_CLK), 				//         hps_io.hps_io_emac1_inst_TX_CLK
        .hps_io_hps_io_emac1_inst_TXD0   (HPS_ENET_TX_DATA[0]),   		//         .hps_io_emac1_inst_TXD0
        .hps_io_hps_io_emac1_inst_TXD1   (HPS_ENET_TX_DATA[1]),   		//         .hps_io_emac1_inst_TXD1
        .hps_io_hps_io_emac1_inst_TXD2   (HPS_ENET_TX_DATA[2]),   		//         .hps_io_emac1_inst_TXD2
        .hps_io_hps_io_emac1_inst_TXD3   (HPS_ENET_TX_DATA[3]),   		//         .hps_io_emac1_inst_TXD3
        .hps_io_hps_io_emac1_inst_RXD0   (HPS_ENET_RX_DATA[0]),   		//         .hps_io_emac1_inst_RXD0
        .hps_io_hps_io_emac1_inst_MDIO   (HPS_ENET_MDIO),   				//         .hps_io_emac1_inst_MDIO
        .hps_io_hps_io_emac1_inst_MDC    (HPS_ENET_MDC),    				//         .hps_io_emac1_inst_MDC
        .hps_io_hps_io_emac1_inst_RX_CTL (HPS_ENET_RX_DV), 					//         .hps_io_emac1_inst_RX_CTL
        .hps_io_hps_io_emac1_inst_TX_CTL (HPS_ENET_TX_EN), 					//         .hps_io_emac1_inst_TX_CTL
        .hps_io_hps_io_emac1_inst_RX_CLK (HPS_ENET_RX_CLK), 				//         .hps_io_emac1_inst_RX_CLK
        .hps_io_hps_io_emac1_inst_RXD1   (HPS_ENET_RX_DATA[1]),   		//         .hps_io_emac1_inst_RXD1
        .hps_io_hps_io_emac1_inst_RXD2   (HPS_ENET_RX_DATA[2]),   		//         .hps_io_emac1_inst_RXD2
        .hps_io_hps_io_emac1_inst_RXD3   (HPS_ENET_RX_DATA[3]),   		//         .hps_io_emac1_inst_RXD3
        .hps_io_hps_io_sdio_inst_CMD     (HPS_SD_CMD),     					//         .hps_io_sdio_inst_CMD
        .hps_io_hps_io_sdio_inst_D0      (HPS_SD_DATA[0]), 			    	//         .hps_io_sdio_inst_D0
        .hps_io_hps_io_sdio_inst_D1      (HPS_SD_DATA[1]),      			//         .hps_io_sdio_inst_D1
        .hps_io_hps_io_sdio_inst_CLK     (HPS_SD_CLK),     					//         .hps_io_sdio_inst_CLK
        .hps_io_hps_io_sdio_inst_D2      (HPS_SD_DATA[2]),    			   //         .hps_io_sdio_inst_D2
        .hps_io_hps_io_sdio_inst_D3      (HPS_SD_DATA[3]),      			//         .hps_io_sdio_inst_D3
        .hps_io_hps_io_usb1_inst_D0      (HPS_USB_DATA[0]),     			//         .hps_io_usb1_inst_D0
        .hps_io_hps_io_usb1_inst_D1      (HPS_USB_DATA[1]),      			//         .hps_io_usb1_inst_D1
        .hps_io_hps_io_usb1_inst_D2      (HPS_USB_DATA[2]),      			//         .hps_io_usb1_inst_D2
        .hps_io_hps_io_usb1_inst_D3      (HPS_USB_DATA[3]),      			//         .hps_io_usb1_inst_D3
        .hps_io_hps_io_usb1_inst_D4      (HPS_USB_DATA[4]),      			//         .hps_io_usb1_inst_D4
        .hps_io_hps_io_usb1_inst_D5      (HPS_USB_DATA[5]),      			//         .hps_io_usb1_inst_D5
        .hps_io_hps_io_usb1_inst_D6      (HPS_USB_DATA[6]),      			//         .hps_io_usb1_inst_D6
        .hps_io_hps_io_usb1_inst_D7      (HPS_USB_DATA[7]),      			//         .hps_io_usb1_inst_D7
        .hps_io_hps_io_usb1_inst_CLK     (HPS_USB_CLKOUT),     			//         .hps_io_usb1_inst_CLK
        .hps_io_hps_io_usb1_inst_STP     (HPS_USB_STP),     				//         .hps_io_usb1_inst_STP
        .hps_io_hps_io_usb1_inst_DIR     (HPS_USB_DIR),     				//         .hps_io_usb1_inst_DIR
        .hps_io_hps_io_usb1_inst_NXT     (HPS_USB_NXT),     				//         .hps_io_usb1_inst_NXT
        .hps_io_hps_io_uart0_inst_RX     (HPS_UART_RX),     				//         .hps_io_uart0_inst_RX
        .hps_io_hps_io_uart0_inst_TX     (HPS_UART_TX),     				//         .hps_io_uart0_inst_TX
        .hps_io_hps_io_gpio_inst_GPIO35  (HPS_ENET_INT_N),  				//         .hps_io_gpio_inst_GPIO35
        .leds_export                     (LEDR),                        //         leds.export
        .memory_0_mem_a                  (HPS_DDR3_ADDR),               //         memory_0.mem_a
        .memory_0_mem_ba                 (HPS_DDR3_BA),                 //         .mem_ba
        .memory_0_mem_ck                 (HPS_DDR3_CK_P),               //         .mem_ck
        .memory_0_mem_ck_n               (HPS_DDR3_CK_N),               //         .mem_ck_n
        .memory_0_mem_cke                (HPS_DDR3_CKE),                //         .mem_cke
        .memory_0_mem_cs_n               (HPS_DDR3_CS_N),               //         .mem_cs_n
        .memory_0_mem_ras_n              (HPS_DDR3_RAS_N),              //         .mem_ras_n
        .memory_0_mem_cas_n              (HPS_DDR3_CAS_N),              //         .mem_cas_n
        .memory_0_mem_we_n               (HPS_DDR3_WE_N),               //         .mem_we_n
        .memory_0_mem_reset_n            (HPS_DDR3_RESET_N),            //         .mem_reset_n
        .memory_0_mem_dq                 (HPS_DDR3_DQ),                 //         .mem_dq
        .memory_0_mem_dqs                (HPS_DDR3_DQS_P),              //         .mem_dqs
        .memory_0_mem_dqs_n              (HPS_DDR3_DQS_N),              //         .mem_dqs_n
        .memory_0_mem_odt                (HPS_DDR3_ODT),                //         .mem_odt
        .memory_0_mem_dm                 (HPS_DDR3_DM),                 //         .mem_dm
        .memory_0_oct_rzqin              (HPS_DDR3_RZQ),                //         .oct_rzqin
        .switches_export                 (SW),                          //         switches.export
        .hex3_export                     (HEX3),                        //         hex3.export
        .hex4_export                     (HEX4),                        //         hex4.export
        .hex5_export                     (HEX5)                         //         hex5.export
    );


	 
endmodule
