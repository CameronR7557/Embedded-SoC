// TermProject.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module TermProject (
		input  wire        clk_clk,                         //     clk.clk
		output wire [6:0]  hex0_export,                     //    hex0.export
		output wire [6:0]  hex1_export,                     //    hex1.export
		output wire [6:0]  hex2_export,                     //    hex2.export
		output wire [6:0]  hex3_export,                     //    hex3.export
		output wire [6:0]  hex4_export,                     //    hex4.export
		output wire [6:0]  hex5_export,                     //    hex5.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //  hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //        .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //        .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //        .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //        .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //        .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //        .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //        .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //        .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //        .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //        .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //        .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //        .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //        .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //        .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //        .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //        .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //        .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //        .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //        .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //        .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //        .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //        .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //        .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //        .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //        .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //        .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //        .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //        .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //        .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //        .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //        .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim0_inst_CLK,    //        .hps_io_spim0_inst_CLK
		output wire        hps_io_hps_io_spim0_inst_MOSI,   //        .hps_io_spim0_inst_MOSI
		input  wire        hps_io_hps_io_spim0_inst_MISO,   //        .hps_io_spim0_inst_MISO
		output wire        hps_io_hps_io_spim0_inst_SS0,    //        .hps_io_spim0_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //        .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //        .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //        .hps_io_gpio_inst_GPIO35
		output wire [14:0] memory_mem_a,                    //  memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //        .mem_ba
		output wire        memory_mem_ck,                   //        .mem_ck
		output wire        memory_mem_ck_n,                 //        .mem_ck_n
		output wire        memory_mem_cke,                  //        .mem_cke
		output wire        memory_mem_cs_n,                 //        .mem_cs_n
		output wire        memory_mem_ras_n,                //        .mem_ras_n
		output wire        memory_mem_cas_n,                //        .mem_cas_n
		output wire        memory_mem_we_n,                 //        .mem_we_n
		output wire        memory_mem_reset_n,              //        .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //        .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //        .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //        .mem_dqs_n
		output wire        memory_mem_odt,                  //        .mem_odt
		output wire [3:0]  memory_mem_dm,                   //        .mem_dm
		input  wire        memory_oct_rzqin,                //        .oct_rzqin
		input  wire        uart_rx_conduit                  // uart_rx.conduit
	);

	wire         clockdivider_0_clock_source_clk;                               // ClockDivider_0:clk_out -> [UART_RX_0:clk, mm_interconnect_0:ClockDivider_0_clock_source_clk, rst_controller_001:clk]
	wire         hps_0_h2f_reset_reset;                                         // hps_0:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                               // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                 // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                 // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                 // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                   // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                               // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                 // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                               // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                               // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                  // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                               // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                 // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                  // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                               // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_clockdivider_0_avalon_slave_0_chipselect;    // mm_interconnect_0:ClockDivider_0_avalon_slave_0_chipselect -> ClockDivider_0:chipselect
	wire   [1:0] mm_interconnect_0_clockdivider_0_avalon_slave_0_address;       // mm_interconnect_0:ClockDivider_0_avalon_slave_0_address -> ClockDivider_0:address
	wire         mm_interconnect_0_clockdivider_0_avalon_slave_0_write;         // mm_interconnect_0:ClockDivider_0_avalon_slave_0_write -> ClockDivider_0:write
	wire  [31:0] mm_interconnect_0_clockdivider_0_avalon_slave_0_writedata;     // mm_interconnect_0:ClockDivider_0_avalon_slave_0_writedata -> ClockDivider_0:writedata
	wire         mm_interconnect_0_uart_rx_0_avalon_slave_0_chipselect;         // mm_interconnect_0:UART_RX_0_avalon_slave_0_chipselect -> UART_RX_0:chipselect
	wire  [31:0] mm_interconnect_0_uart_rx_0_avalon_slave_0_readdata;           // UART_RX_0:readdata -> mm_interconnect_0:UART_RX_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_uart_rx_0_avalon_slave_0_address;            // mm_interconnect_0:UART_RX_0_avalon_slave_0_address -> UART_RX_0:address
	wire         mm_interconnect_0_uart_rx_0_avalon_slave_0_read;               // mm_interconnect_0:UART_RX_0_avalon_slave_0_read -> UART_RX_0:read
	wire         mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_chipselect -> SevenSegDecoder_4:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_address -> SevenSegDecoder_4:address
	wire         mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_write -> SevenSegDecoder_4:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_4_avalon_slave_0_writedata -> SevenSegDecoder_4:writedata
	wire         mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_chipselect -> SevenSegDecoder_3:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_address -> SevenSegDecoder_3:address
	wire         mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_write -> SevenSegDecoder_3:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_3_avalon_slave_0_writedata -> SevenSegDecoder_3:writedata
	wire         mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_chipselect -> SevenSegDecoder_2:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_address -> SevenSegDecoder_2:address
	wire         mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_write -> SevenSegDecoder_2:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_2_avalon_slave_0_writedata -> SevenSegDecoder_2:writedata
	wire         mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_chipselect -> SevenSegDecoder_1:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_address -> SevenSegDecoder_1:address
	wire         mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_write -> SevenSegDecoder_1:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_1_avalon_slave_0_writedata -> SevenSegDecoder_1:writedata
	wire         mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_chipselect -> SevenSegDecoder_0:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_address -> SevenSegDecoder_0:address
	wire         mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_write -> SevenSegDecoder_0:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_0_avalon_slave_0_writedata -> SevenSegDecoder_0:writedata
	wire         mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect; // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_chipselect -> SevenSegDecoder_5:chipselect
	wire   [1:0] mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address;    // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_address -> SevenSegDecoder_5:address
	wire         mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write;      // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_write -> SevenSegDecoder_5:write
	wire  [31:0] mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata;  // mm_interconnect_0:SevenSegDecoder_5_avalon_slave_0_writedata -> SevenSegDecoder_5:writedata
	wire         mm_interconnect_0_crc_0_avalon_slave_0_chipselect;             // mm_interconnect_0:CRC_0_avalon_slave_0_chipselect -> CRC_0:chipselect
	wire  [31:0] mm_interconnect_0_crc_0_avalon_slave_0_readdata;               // CRC_0:readdata -> mm_interconnect_0:CRC_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_crc_0_avalon_slave_0_address;                // mm_interconnect_0:CRC_0_avalon_slave_0_address -> CRC_0:address
	wire         mm_interconnect_0_crc_0_avalon_slave_0_read;                   // mm_interconnect_0:CRC_0_avalon_slave_0_read -> CRC_0:read
	wire         mm_interconnect_0_crc_0_avalon_slave_0_write;                  // mm_interconnect_0:CRC_0_avalon_slave_0_write -> CRC_0:write
	wire  [31:0] mm_interconnect_0_crc_0_avalon_slave_0_writedata;              // mm_interconnect_0:CRC_0_avalon_slave_0_writedata -> CRC_0:writedata
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [CRC_0:reset_n, ClockDivider_0:reset_n, SevenSegDecoder_0:reset_n, SevenSegDecoder_1:reset_n, SevenSegDecoder_2:reset_n, SevenSegDecoder_3:reset_n, SevenSegDecoder_4:reset_n, SevenSegDecoder_5:reset_n, mm_interconnect_0:ClockDivider_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [UART_RX_0:reset_n, mm_interconnect_0:UART_RX_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	My_CRC crc_0 (
		.clk        (clk_clk),                                           //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.address    (mm_interconnect_0_crc_0_avalon_slave_0_address),    // avalon_slave_0.address
		.read       (mm_interconnect_0_crc_0_avalon_slave_0_read),       //               .read
		.write      (mm_interconnect_0_crc_0_avalon_slave_0_write),      //               .write
		.chipselect (mm_interconnect_0_crc_0_avalon_slave_0_chipselect), //               .chipselect
		.writedata  (mm_interconnect_0_crc_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_crc_0_avalon_slave_0_readdata)    //               .readdata
	);

	My_ClockDivider clockdivider_0 (
		.clk        (clk_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //          reset.reset_n
		.chipselect (mm_interconnect_0_clockdivider_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.address    (mm_interconnect_0_clockdivider_0_avalon_slave_0_address),    //               .address
		.write      (mm_interconnect_0_clockdivider_0_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_clockdivider_0_avalon_slave_0_writedata),  //               .writedata
		.clk_out    (clockdivider_0_clock_source_clk)                             //   clock_source.clk
	);

	SevenSegDecoder sevensegdecoder_0 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex0_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_1 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex1_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_2 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex2_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_3 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex3_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_4 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex4_export)                                                    //    conduit_end.export
	);

	SevenSegDecoder sevensegdecoder_5 (
		.clk        (clk_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                               //          reset.reset_n
		.address    (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address),    // avalon_slave_0.address
		.write      (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata),  //               .writedata
		.chipselect (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect), //               .chipselect
		.segs       (hex5_export)                                                    //    conduit_end.export
	);

	My_UART_RX uart_rx_0 (
		.clk        (clockdivider_0_clock_source_clk),                       //          clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //          reset.reset_n
		.address    (mm_interconnect_0_uart_rx_0_avalon_slave_0_address),    // avalon_slave_0.address
		.read       (mm_interconnect_0_uart_rx_0_avalon_slave_0_read),       //               .read
		.chipselect (mm_interconnect_0_uart_rx_0_avalon_slave_0_chipselect), //               .chipselect
		.readdata   (mm_interconnect_0_uart_rx_0_avalon_slave_0_readdata),   //               .readdata
		.RX_in      (uart_rx_conduit)                                        //    conduit_end.conduit
	);

	TermProject_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_io_hps_io_spim0_inst_CLK),    //                  .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_io_hps_io_spim0_inst_MOSI),   //                  .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_io_hps_io_spim0_inst_MISO),   //                  .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_io_hps_io_spim0_inst_SS0),    //                  .hps_io_spim0_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	TermProject_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                  //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                 //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                               //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                               //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                               //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                               //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                   //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                 //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                 //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                 //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                   //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                 //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                  //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                 //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                               //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                               //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                               //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                               //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                   //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                 //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                 //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                 //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                       //                                                     clk_0_clk.clk
		.ClockDivider_0_clock_source_clk                                     (clockdivider_0_clock_source_clk),                               //                                   ClockDivider_0_clock_source.clk
		.ClockDivider_0_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                                //                    ClockDivider_0_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                            // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.UART_RX_0_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                            //                         UART_RX_0_reset_reset_bridge_in_reset.reset
		.ClockDivider_0_avalon_slave_0_address                               (mm_interconnect_0_clockdivider_0_avalon_slave_0_address),       //                                 ClockDivider_0_avalon_slave_0.address
		.ClockDivider_0_avalon_slave_0_write                                 (mm_interconnect_0_clockdivider_0_avalon_slave_0_write),         //                                                              .write
		.ClockDivider_0_avalon_slave_0_writedata                             (mm_interconnect_0_clockdivider_0_avalon_slave_0_writedata),     //                                                              .writedata
		.ClockDivider_0_avalon_slave_0_chipselect                            (mm_interconnect_0_clockdivider_0_avalon_slave_0_chipselect),    //                                                              .chipselect
		.CRC_0_avalon_slave_0_address                                        (mm_interconnect_0_crc_0_avalon_slave_0_address),                //                                          CRC_0_avalon_slave_0.address
		.CRC_0_avalon_slave_0_write                                          (mm_interconnect_0_crc_0_avalon_slave_0_write),                  //                                                              .write
		.CRC_0_avalon_slave_0_read                                           (mm_interconnect_0_crc_0_avalon_slave_0_read),                   //                                                              .read
		.CRC_0_avalon_slave_0_readdata                                       (mm_interconnect_0_crc_0_avalon_slave_0_readdata),               //                                                              .readdata
		.CRC_0_avalon_slave_0_writedata                                      (mm_interconnect_0_crc_0_avalon_slave_0_writedata),              //                                                              .writedata
		.CRC_0_avalon_slave_0_chipselect                                     (mm_interconnect_0_crc_0_avalon_slave_0_chipselect),             //                                                              .chipselect
		.SevenSegDecoder_0_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_address),    //                              SevenSegDecoder_0_avalon_slave_0.address
		.SevenSegDecoder_0_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_0_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_0_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_0_avalon_slave_0_chipselect), //                                                              .chipselect
		.SevenSegDecoder_1_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_address),    //                              SevenSegDecoder_1_avalon_slave_0.address
		.SevenSegDecoder_1_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_1_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_1_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_1_avalon_slave_0_chipselect), //                                                              .chipselect
		.SevenSegDecoder_2_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_address),    //                              SevenSegDecoder_2_avalon_slave_0.address
		.SevenSegDecoder_2_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_2_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_2_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_2_avalon_slave_0_chipselect), //                                                              .chipselect
		.SevenSegDecoder_3_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_address),    //                              SevenSegDecoder_3_avalon_slave_0.address
		.SevenSegDecoder_3_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_3_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_3_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_3_avalon_slave_0_chipselect), //                                                              .chipselect
		.SevenSegDecoder_4_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_address),    //                              SevenSegDecoder_4_avalon_slave_0.address
		.SevenSegDecoder_4_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_4_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_4_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_4_avalon_slave_0_chipselect), //                                                              .chipselect
		.SevenSegDecoder_5_avalon_slave_0_address                            (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_address),    //                              SevenSegDecoder_5_avalon_slave_0.address
		.SevenSegDecoder_5_avalon_slave_0_write                              (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_write),      //                                                              .write
		.SevenSegDecoder_5_avalon_slave_0_writedata                          (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_writedata),  //                                                              .writedata
		.SevenSegDecoder_5_avalon_slave_0_chipselect                         (mm_interconnect_0_sevensegdecoder_5_avalon_slave_0_chipselect), //                                                              .chipselect
		.UART_RX_0_avalon_slave_0_address                                    (mm_interconnect_0_uart_rx_0_avalon_slave_0_address),            //                                      UART_RX_0_avalon_slave_0.address
		.UART_RX_0_avalon_slave_0_read                                       (mm_interconnect_0_uart_rx_0_avalon_slave_0_read),               //                                                              .read
		.UART_RX_0_avalon_slave_0_readdata                                   (mm_interconnect_0_uart_rx_0_avalon_slave_0_readdata),           //                                                              .readdata
		.UART_RX_0_avalon_slave_0_chipselect                                 (mm_interconnect_0_uart_rx_0_avalon_slave_0_chipselect)          //                                                              .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clockdivider_0_clock_source_clk),    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
