// Lab04.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module Lab04 (
		input  wire        clk_clk,            //         clk.clk
		output wire [9:0]  leds_export,        //        leds.export
		input  wire [3:0]  pushbuttons_export, // pushbuttons.export
		output wire        sdram_clk_clk,      //   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,    //  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,      //            .ba
		output wire        sdram_wire_cas_n,   //            .cas_n
		output wire        sdram_wire_cke,     //            .cke
		output wire        sdram_wire_cs_n,    //            .cs_n
		inout  wire [15:0] sdram_wire_dq,      //            .dq
		output wire [1:0]  sdram_wire_dqm,     //            .dqm
		output wire        sdram_wire_ras_n,   //            .ras_n
		output wire        sdram_wire_we_n     //            .we_n
	);

	wire         clocks_sys_clk_clk;                                    // CLOCKS:sys_clk_clk -> [DEBUG:clk, LEDs:clk, Lab04:clk, SDRAM:clk, irq_mapper:clk, mm_interconnect_0:CLOCKS_sys_clk_clk, pushbuttons:clk, rst_controller:clk, sys_clk:clk]
	wire         lab04_debug_reset_request_reset;                       // Lab04:debug_reset_request -> [CLOCKS:ref_reset_reset, rst_controller:reset_in0]
	wire  [31:0] lab04_data_master_readdata;                            // mm_interconnect_0:Lab04_data_master_readdata -> Lab04:d_readdata
	wire         lab04_data_master_waitrequest;                         // mm_interconnect_0:Lab04_data_master_waitrequest -> Lab04:d_waitrequest
	wire         lab04_data_master_debugaccess;                         // Lab04:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Lab04_data_master_debugaccess
	wire  [27:0] lab04_data_master_address;                             // Lab04:d_address -> mm_interconnect_0:Lab04_data_master_address
	wire   [3:0] lab04_data_master_byteenable;                          // Lab04:d_byteenable -> mm_interconnect_0:Lab04_data_master_byteenable
	wire         lab04_data_master_read;                                // Lab04:d_read -> mm_interconnect_0:Lab04_data_master_read
	wire         lab04_data_master_write;                               // Lab04:d_write -> mm_interconnect_0:Lab04_data_master_write
	wire  [31:0] lab04_data_master_writedata;                           // Lab04:d_writedata -> mm_interconnect_0:Lab04_data_master_writedata
	wire  [31:0] lab04_instruction_master_readdata;                     // mm_interconnect_0:Lab04_instruction_master_readdata -> Lab04:i_readdata
	wire         lab04_instruction_master_waitrequest;                  // mm_interconnect_0:Lab04_instruction_master_waitrequest -> Lab04:i_waitrequest
	wire  [27:0] lab04_instruction_master_address;                      // Lab04:i_address -> mm_interconnect_0:Lab04_instruction_master_address
	wire         lab04_instruction_master_read;                         // Lab04:i_read -> mm_interconnect_0:Lab04_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_lab04_debug_mem_slave_readdata;      // Lab04:debug_mem_slave_readdata -> mm_interconnect_0:Lab04_debug_mem_slave_readdata
	wire         mm_interconnect_0_lab04_debug_mem_slave_waitrequest;   // Lab04:debug_mem_slave_waitrequest -> mm_interconnect_0:Lab04_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_lab04_debug_mem_slave_debugaccess;   // mm_interconnect_0:Lab04_debug_mem_slave_debugaccess -> Lab04:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_lab04_debug_mem_slave_address;       // mm_interconnect_0:Lab04_debug_mem_slave_address -> Lab04:debug_mem_slave_address
	wire         mm_interconnect_0_lab04_debug_mem_slave_read;          // mm_interconnect_0:Lab04_debug_mem_slave_read -> Lab04:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_lab04_debug_mem_slave_byteenable;    // mm_interconnect_0:Lab04_debug_mem_slave_byteenable -> Lab04:debug_mem_slave_byteenable
	wire         mm_interconnect_0_lab04_debug_mem_slave_write;         // mm_interconnect_0:Lab04_debug_mem_slave_write -> Lab04:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_lab04_debug_mem_slave_writedata;     // mm_interconnect_0:Lab04_debug_mem_slave_writedata -> Lab04:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                 // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                   // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                    // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                       // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                 // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;              // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                      // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                  // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_sys_clk_s1_chipselect;               // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                 // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                  // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                    // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                  // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                    // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [2:0] mm_interconnect_0_leds_s1_address;                     // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                       // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                   // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;             // pushbuttons:readdata -> mm_interconnect_0:pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;              // mm_interconnect_0:pushbuttons_s1_address -> pushbuttons:address
	wire         irq_mapper_receiver0_irq;                              // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                              // sys_clk:irq -> irq_mapper:receiver1_irq
	wire  [31:0] lab04_irq_irq;                                         // irq_mapper:sender_irq -> Lab04:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [DEBUG:rst_n, LEDs:reset_n, Lab04:reset_n, SDRAM:reset_n, irq_mapper:reset, mm_interconnect_0:Lab04_reset_reset_bridge_in_reset_reset, pushbuttons:reset_n, rst_translator:in_reset, sys_clk:reset_n]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [Lab04:reset_req, rst_translator:reset_req_in]

	Lab04_CLOCKS clocks (
		.ref_clk_clk        (clk_clk),                         //      ref_clk.clk
		.ref_reset_reset    (lab04_debug_reset_request_reset), //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),              //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                   //    sdram_clk.clk
		.reset_source_reset ()                                 // reset_source.reset
	);

	Lab04_DEBUG debug (
		.clk            (clocks_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	Lab04_LEDs leds (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	Lab04_Lab04 lab04 (
		.clk                                 (clocks_sys_clk_clk),                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (lab04_data_master_address),                           //               data_master.address
		.d_byteenable                        (lab04_data_master_byteenable),                        //                          .byteenable
		.d_read                              (lab04_data_master_read),                              //                          .read
		.d_readdata                          (lab04_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (lab04_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (lab04_data_master_write),                             //                          .write
		.d_writedata                         (lab04_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (lab04_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (lab04_instruction_master_address),                    //        instruction_master.address
		.i_read                              (lab04_instruction_master_read),                       //                          .read
		.i_readdata                          (lab04_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (lab04_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (lab04_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (lab04_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_lab04_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_lab04_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_lab04_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_lab04_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_lab04_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_lab04_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_lab04_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_lab04_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	Lab04_SDRAM sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Lab04_pushbuttons pushbuttons (
		.clk      (clocks_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pushbuttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pushbuttons_s1_readdata), //                    .readdata
		.in_port  (pushbuttons_export)                         // external_connection.export
	);

	Lab04_sys_clk sys_clk (
		.clk        (clocks_sys_clk_clk),                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	Lab04_mm_interconnect_0 mm_interconnect_0 (
		.CLOCKS_sys_clk_clk                      (clocks_sys_clk_clk),                                    //                    CLOCKS_sys_clk.clk
		.Lab04_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // Lab04_reset_reset_bridge_in_reset.reset
		.Lab04_data_master_address               (lab04_data_master_address),                             //                 Lab04_data_master.address
		.Lab04_data_master_waitrequest           (lab04_data_master_waitrequest),                         //                                  .waitrequest
		.Lab04_data_master_byteenable            (lab04_data_master_byteenable),                          //                                  .byteenable
		.Lab04_data_master_read                  (lab04_data_master_read),                                //                                  .read
		.Lab04_data_master_readdata              (lab04_data_master_readdata),                            //                                  .readdata
		.Lab04_data_master_write                 (lab04_data_master_write),                               //                                  .write
		.Lab04_data_master_writedata             (lab04_data_master_writedata),                           //                                  .writedata
		.Lab04_data_master_debugaccess           (lab04_data_master_debugaccess),                         //                                  .debugaccess
		.Lab04_instruction_master_address        (lab04_instruction_master_address),                      //          Lab04_instruction_master.address
		.Lab04_instruction_master_waitrequest    (lab04_instruction_master_waitrequest),                  //                                  .waitrequest
		.Lab04_instruction_master_read           (lab04_instruction_master_read),                         //                                  .read
		.Lab04_instruction_master_readdata       (lab04_instruction_master_readdata),                     //                                  .readdata
		.DEBUG_avalon_jtag_slave_address         (mm_interconnect_0_debug_avalon_jtag_slave_address),     //           DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write           (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                  .write
		.DEBUG_avalon_jtag_slave_read            (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                  .read
		.DEBUG_avalon_jtag_slave_readdata        (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                  .readdata
		.DEBUG_avalon_jtag_slave_writedata       (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                  .writedata
		.DEBUG_avalon_jtag_slave_waitrequest     (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect      (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.Lab04_debug_mem_slave_address           (mm_interconnect_0_lab04_debug_mem_slave_address),       //             Lab04_debug_mem_slave.address
		.Lab04_debug_mem_slave_write             (mm_interconnect_0_lab04_debug_mem_slave_write),         //                                  .write
		.Lab04_debug_mem_slave_read              (mm_interconnect_0_lab04_debug_mem_slave_read),          //                                  .read
		.Lab04_debug_mem_slave_readdata          (mm_interconnect_0_lab04_debug_mem_slave_readdata),      //                                  .readdata
		.Lab04_debug_mem_slave_writedata         (mm_interconnect_0_lab04_debug_mem_slave_writedata),     //                                  .writedata
		.Lab04_debug_mem_slave_byteenable        (mm_interconnect_0_lab04_debug_mem_slave_byteenable),    //                                  .byteenable
		.Lab04_debug_mem_slave_waitrequest       (mm_interconnect_0_lab04_debug_mem_slave_waitrequest),   //                                  .waitrequest
		.Lab04_debug_mem_slave_debugaccess       (mm_interconnect_0_lab04_debug_mem_slave_debugaccess),   //                                  .debugaccess
		.LEDs_s1_address                         (mm_interconnect_0_leds_s1_address),                     //                           LEDs_s1.address
		.LEDs_s1_write                           (mm_interconnect_0_leds_s1_write),                       //                                  .write
		.LEDs_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                    //                                  .readdata
		.LEDs_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                   //                                  .writedata
		.LEDs_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                  //                                  .chipselect
		.pushbuttons_s1_address                  (mm_interconnect_0_pushbuttons_s1_address),              //                    pushbuttons_s1.address
		.pushbuttons_s1_readdata                 (mm_interconnect_0_pushbuttons_s1_readdata),             //                                  .readdata
		.SDRAM_s1_address                        (mm_interconnect_0_sdram_s1_address),                    //                          SDRAM_s1.address
		.SDRAM_s1_write                          (mm_interconnect_0_sdram_s1_write),                      //                                  .write
		.SDRAM_s1_read                           (mm_interconnect_0_sdram_s1_read),                       //                                  .read
		.SDRAM_s1_readdata                       (mm_interconnect_0_sdram_s1_readdata),                   //                                  .readdata
		.SDRAM_s1_writedata                      (mm_interconnect_0_sdram_s1_writedata),                  //                                  .writedata
		.SDRAM_s1_byteenable                     (mm_interconnect_0_sdram_s1_byteenable),                 //                                  .byteenable
		.SDRAM_s1_readdatavalid                  (mm_interconnect_0_sdram_s1_readdatavalid),              //                                  .readdatavalid
		.SDRAM_s1_waitrequest                    (mm_interconnect_0_sdram_s1_waitrequest),                //                                  .waitrequest
		.SDRAM_s1_chipselect                     (mm_interconnect_0_sdram_s1_chipselect),                 //                                  .chipselect
		.sys_clk_s1_address                      (mm_interconnect_0_sys_clk_s1_address),                  //                        sys_clk_s1.address
		.sys_clk_s1_write                        (mm_interconnect_0_sys_clk_s1_write),                    //                                  .write
		.sys_clk_s1_readdata                     (mm_interconnect_0_sys_clk_s1_readdata),                 //                                  .readdata
		.sys_clk_s1_writedata                    (mm_interconnect_0_sys_clk_s1_writedata),                //                                  .writedata
		.sys_clk_s1_chipselect                   (mm_interconnect_0_sys_clk_s1_chipselect)                //                                  .chipselect
	);

	Lab04_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (lab04_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (lab04_debug_reset_request_reset),    // reset_in0.reset
		.clk            (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
